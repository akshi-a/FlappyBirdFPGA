module LFSR6_testbench();
  
  reg reset, clk; 
  wire [5:0]number;
  
  LFSR6 ch (clk,reset,number);

  // Set up the clock
  parameter CLOCK_PERIOD=100;
  initial clk=1;
  always begin
    #(CLOCK_PERIOD/2); clk = ~clk;
  end
  // Set up the inputs to the design (each line is a clock cycle)
  initial begin
	 @(posedge clk); reset<=1;
	 @(posedge clk); reset<=0;
    for(int i =0; i<64 ; i++) @(posedge clk);
	 @(posedge clk); 
	 @(posedge clk);
	 @(posedge clk);reset<=1;
	 @(posedge clk);reset<=0;
	 @(posedge clk);
	 @(posedge clk);
	 $stop;       // End the simulation
  end 
  
endmodule 